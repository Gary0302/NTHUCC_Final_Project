`timescale 1ns/1ps
module ALU
(
    input [7:0] A,
    input [7:0] B,
    input [3:0] instruction,
    output reg [7:0] F
);
    //TODO: write your design below

endmodule